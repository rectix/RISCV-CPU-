`timescale 1ns / 1ps




`define XLEN          32                 
`define ILEN          32   
`define PC_INIT       32'h0000_0000  
`define NOP_INSTRUCT  32'h0000_0000          


`define XLSB          $clog2(`XLEN/8)-1:0 
